`include "seq_item.sv"
`include "sequence.sv"
`include "seq_full_rw.sv"
`include "seq_7bit.sv"
`include "seq_10bit.sv"
`include "seq_rpt_start.sv"
`include "seq_mismatch.sv"
`include "seq_data_override.sv"
`include "seq_directed.sv"
`include "stuck.sv"

`include "seq_coverpoint.sv"
`include "seq_covercross.sv"
`include "seq_covergroup.sv"
`include "sequencer.sv"
`include "driver.sv"
`include "monitor.sv"
`include "agent.sv"
`include "scoreboard.sv"
`include "coverage.sv"
`include "environment.sv"
`include "test.sv"
