`include "seq_item.sv"
`include "seq_item1.sv"
`include "sequence.sv"
`include "sequence1.sv"
`include "seq_full_rw.sv"
`include "seq_7bit.sv"
`include "seq_10bit.sv"
`include "seq_rpt_start.sv"
`include "seq_mismatch.sv"
`include "seq_data_override.sv"
`include "seq_directed.sv"
`include "stuck.sv"

`include "seq_coverpoint.sv"
`include "seq_covercross.sv"
`include "seq_covergroup.sv"
`include "seq_coverpoint1.sv"
`include "seq_covercross1.sv"
`include "seq_covergroup1.sv"
`include "seq_covercross2.sv"
`include "seq_covergroup2.sv"

`include "sequencer.sv"
`include "driver.sv"
`include "monitor.sv"
`include "agent.sv"
`include "scoreboard.sv"
`include "coverage.sv"
`include "sequencer1.sv"
`include "driver1.sv"
`include "monitor1.sv"
`include "agent1.sv"
`include "scoreboard1.sv"
`include "coverage1.sv"
`include "environment.sv"
`include "test.sv"
